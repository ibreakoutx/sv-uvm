`include "tb_env.sv"
