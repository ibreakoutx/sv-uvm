`define RAL_TB_ENV tb_env

`include "tb_env.sv"
